//Verilog HDL for "comparator", "comp" "functional"


module comp ( vout, \v+ , \v- , vdd, vss );

  input \v+ ;
  output vout;
  input \v- ;
  input vdd;
  input vss;
endmodule
